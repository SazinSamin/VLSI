module sb(su
