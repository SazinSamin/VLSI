module pattern(o, i, rst, clk);
	output reg o;
	input i, rst, clk;
	reg[1:0] states;
	
	 
