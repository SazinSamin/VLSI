module vector;
	reg [7:0] arr[7:0]; // have 8 arr (arr[0], arr[1], ... arr[7]), each 8 bit long
	arr[1] = 34234;

endmodule
