module decoder(out, in, en);
	input in, en;
	output[
