module Parameter;
	parameter N = 4;
	reg out[N-1:0];
	
endmodule
