module exorGate(
			input		a_i,
			input		b_i,
			output		c_o
);

assign c_o = a_i ^ b_i;

endmodule
