module string;
	initial begin
		$display("Verilog is good for learning");
		$display("SystemVerilog is good for testing");
	end
endmodule
