module structure;
	//  defination of structure
	typedef struct {
		int taka;
		real poisa;
	} money;
	
	//  declearation of a structure variable
	money moneyBag;
	
	moneyBag = '{10, 12};
	
endmodule
	
